library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rra_servo_controller is
  generic(
      STEP    : integer
    );
  port(
      i_clk   : in  std_ulogic;
      i_rst   : in  std_ulogic;

      i_speed   	: in  std_ulogic_vector(3 downto 0);
		i_offset 	: in std_ulogic_vector(7 downto 0);
      o_current 	: out std_ulogic_vector(9 downto 0);
	   o_current_i	: out std_ulogic_vector(9 downto 0);
      i_target  	: in  std_ulogic_vector(9 downto 0);
      o_pwm_out 	: out std_ulogic;
	   o_pwm_out_i	: out std_ulogic
    );
  
end rra_servo_controller;

architecture rtl of rra_servo_controller is
  signal current: integer range 0 to 2000;
  signal current_i : integer range 0 to 2000;
  signal target: integer range 0 to 2000;
  signal speed: unsigned(3 downto 0);
  signal pwm_out:   std_ulogic;
  signal pwm_out_i:   std_ulogic;

  signal interval: integer range 0 to 2000;
  signal interval_count: integer range 0 to 2000;

  signal pwm_count: integer range 0 to 20000;
  signal pwm_count_i: integer range 0 to 20000;

  signal clk_1mhz: std_ulogic;
  signal clk_1khz: std_ulogic;
  signal clk_1mhz_count: integer range 0 to 49;
  signal clk_1khz_count: integer range 0 to 999;

begin

  move: process(i_rst, clk_1khz)
  begin
    if i_rst = '1' then
      current <= 0;
      target <= 0;
      speed <= (others => '0');

      o_current <= (others => '0');

      interval_count <= 0;
      interval <= 991;
    else
      if rising_edge(clk_1khz) then

          interval <= (((to_integer(unsigned(i_speed)) * 62) + 62) - 1);

          if interval_count < interval then
            interval_count <= interval_count + 1;
          else
            if current = target then
              --Do nothing
            elsif current < target then
              --Check to see if increment would jump over target
              if (current + STEP) > target then
                --If it does, assign the target (partial step)
                current <= target;
              else
                --If not, increment by the full step
                --current <= current + STEP;
					 current <= target;
              end if;
            elsif current > target then
              --Check to see if decrement would jump over target
              if (current - STEP) < target then
                --If it does, assign the target (partial step)
                current <= target;
              else
                --If not, decrement by the full step
                --current <= current - STEP;
					 current <= target;
              end if;
            end if;
            interval_count <= 0;
          end if;
        end if;

        speed <= unsigned(i_speed);
        target <= to_integer(unsigned(i_target));
        o_current <= std_ulogic_vector(to_unsigned(current, o_current'length));
		o_current_i <= std_ulogic_vector(to_unsigned(current_i, o_current_i'length));
      end if;
  end process;


  clocks: process(i_clk)  
  begin
    if rising_edge(i_clk) then
      if i_rst = '1' then
        clk_1mhz_count <= 0;
        clk_1mhz <= '0';
        clk_1khz_count <= 0;
        clk_1khz <= '0';
      else
      --1mhz clock
        if clk_1mhz_count < 49 then
          clk_1mhz_count <= clk_1mhz_count + 1;
          clk_1mhz <= '0';
        else
          clk_1mhz_count <= 0;
          clk_1mhz <= '1';

          --1kHz clock
          if clk_1khz_count < 999 then
            clk_1khz_count <= clk_1khz_count + 1;
            clk_1khz <= '0';
          else  
            clk_1khz_count <= 0;
            clk_1khz <= '1';
          end if;
        end if;
      end if;
    end if;
  end process;

  pwm: process(i_clk, clk_1mhz)
  begin

    if i_rst = '1' then
      pwm_out <= '0';
      o_pwm_out <= '0';
      pwm_count <= 0;
    else
      if rising_edge(clk_1mhz) then
        if pwm_count < 1000 then
          --Stay high for at least 1ms
          pwm_count <= pwm_count + 1;
          pwm_out <= '1';
        elsif pwm_count < (1000 + (current)) then
          pwm_count <= pwm_count + 1;
          pwm_out <= '1';
        elsif pwm_count < 20000 then
          pwm_count <= pwm_count + 1;
          pwm_out <= '0';
        else
          pwm_count <= 0;
          pwm_out <= '0';
        end if;
      end if;

      if rising_edge(i_clk) then
        o_pwm_out <= pwm_out;
      end if;
    end if;
  end process;
  
  pwm_i: process(i_clk, clk_1mhz)
  begin

    if i_rst = '1' then
      pwm_out_i <= '0';
      o_pwm_out_i <= '0';
      pwm_count_i <= 0;
    else
      if rising_edge(clk_1mhz) then
        if pwm_count_i < 1000 then
          --Stay high for at least 1ms
          pwm_count_i <= pwm_count_i + 1;
          pwm_out_i <= '1';
        elsif pwm_count_i < (1000 + current_i + (to_integer(signed(i_offset)))) then
          pwm_count_i <= pwm_count_i + 1;
          pwm_out_i <= '1';
        elsif pwm_count_i < 20000 then
          pwm_count_i <= pwm_count_i + 1;
          pwm_out_i <= '0';
        else
          pwm_count_i <= 0;
          pwm_out_i <= '0';
        end if;
      end if;

      if rising_edge(i_clk) then
        o_pwm_out_i <= pwm_out_i;
      end if;
    end if;
  end process;
  
  current_i <= 991 - current;
end rtl;

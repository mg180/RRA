library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity rra is
port (
		clk			: in  std_ulogic;
		rst			: in  std_ulogic;

		--Servo Positions
		l1,l2		: out std_ulogic;	
		m1,m2		: out std_ulogic;
		u1,u2		: out std_ulogic;
		w1,g1 	: out std_ulogic;
		b1			: out std_ulogic;

		--Control
		low_u		: in std_ulogic;
		low_d		: in std_ulogic;
		mid_u		: in std_ulogic;
		mid_d		: in std_ulogic;
		upp_u		: in std_ulogic;
		upp_d		: in std_ulogic;
		store 		: in std_ulogic;
	   low_target : out std_logic_vector(8 downto 0);
		speed		: in std_ulogic_vector(3 downto 0);
		mode		: in std_ulogic_vector(1 downto 0)
	 );
end rra;

architecture v1 of rra is

	component rra_memory
	port(
			clk		: in  std_ulogic;
			rst 	: in  std_ulogic;

			addr	: in  std_ulogic_vector(7 downto 0);
			data_in	: in  std_ulogic_vector(63 downto 0);
			data_out: out std_ulogic_vector(63 downto 0);
			l_memory: in  std_ulogic;
			w_memory: in  std_ulogic
		);
	end component;

	component controller
	port(
			clk       : in  std_ulogic;
	        rst       : in  std_ulogic;
	        
	        mode      : in  std_ulogic_vector(1 downto 0);
	        moving    : in  std_ulogic;
	        store     : in  std_ulogic;
	        l_keypad  : out std_ulogic;
	        l_memory  : out std_ulogic;
	        w_memory  : out std_ulogic
		);
	end component;

	component rra_servo_controller
	generic(
			STEP		: integer
		);
	port(
			i_clk		: in  std_ulogic;
			i_rst		: in  std_ulogic;

			i_speed 	: in  std_ulogic_vector(3 downto 0);
			o_current	: out unsigned(8 downto 0);
			i_target  	: in  unsigned(8 downto 0);
			o_pwm_out 	: out std_ulogic
		);
	end component;

	--Memory
	signal addr		: std_ulogic_vector(7 downto 0);
	signal data_in	: std_ulogic_vector(63 downto 0);
	signal data_out	: std_ulogic_vector(63 downto 0);
	signal l_memory : std_ulogic;
	signal w_memory : std_ulogic;

	--Movement (c - current, t - target)
	constant SERVO_STEP					: integer := 10;
	signal moving						: std_ulogic;
	signal c_lower_pos,		t_lower_pos	: unsigned(8 downto 0);
	signal c_middle_pos,	t_middle_pos: unsigned(8 downto 0);
	signal c_upper_pos,		t_upper_pos	: unsigned(8 downto 0);
	signal c_wrist_pos,		t_wrist_pos	: unsigned(8 downto 0);
	signal c_gripper_pos,		t_gripper_pos	: unsigned(8 downto 0);
	signal c_base_pos,		t_base_pos	: unsigned(8 downto 0);

	--Servo control
	signal l_keypad 					: std_ulogic;
	signal l_pwm, m_pwm, u_pwm, g_pwm, b_pwm, w_pwm			: std_ulogic;

begin
	
	memory : rra_memory	 
	port map(
		clk 		=> clk,
		rst 		=> rst,
		addr		=> addr,
		data_in		=> data_in,
		data_out	=> data_out,
		l_memory	=> l_memory,
		w_memory	=> w_memory
	);

	rra_controller	: controller 
	port map(
		clk 		=> clk,
		rst 		=> rst,
		mode 		=> mode,
		moving  	=> moving,
		store 		=> store,
		l_keypad	=> l_keypad,
		l_memory	=> l_memory,
		w_memory	=> w_memory
	);

	rra_servo_lower : rra_servo_controller 
	generic map(
		STEP 		=> SERVO_STEP
	)
	port map(
		i_clk 		=> clk,
		i_rst 		=> rst,
		i_speed		=> speed,
		o_current	=> c_lower_pos,
		i_target	=> t_lower_pos,
		o_pwm_out	=> l_pwm
	);

	rra_servo_middle: rra_servo_controller 
	generic map(
		STEP 		=> SERVO_STEP
	)
	port map(
		i_clk 		=> clk,
		i_rst 		=> rst,
		i_speed		=> speed,
		o_current	=> c_lower_pos,
		i_target	=> t_lower_pos,
		o_pwm_out	=> m_pwm
	);

	rra_servo_upper : rra_servo_controller 
	generic map(
		STEP 		=> SERVO_STEP
	)
	port map(
		i_clk 		=> clk,
		i_rst 		=> rst,
		i_speed		=> speed,
		o_current	=> c_lower_pos,
		i_target	=> t_lower_pos,
		o_pwm_out	=> u_pwm
	);
	
   rra_servo_wrist : rra_servo_controller 
	generic map(
		STEP 		=> SERVO_STEP
	)
	port map(
		i_clk 		=> clk,
		i_rst 		=> rst,
		i_speed		=> speed,
		o_current	=> c_wrist_pos,
		i_target	=> t_wrist_pos,
		o_pwm_out	=> w_pwm
	);
	
	rra_servo_gripper : rra_servo_controller 
	generic map(
		STEP 		=> SERVO_STEP
	)
	port map(
		i_clk 		=> clk,
		i_rst 		=> rst,
		i_speed		=> speed,
		o_current	=> c_gripper_pos,
		i_target	=> t_gripper_pos,
		o_pwm_out	=> g_pwm
	);
	
	rra_servo_base : rra_servo_controller 
	generic map(
		STEP 		=> SERVO_STEP
	)
	port map(
		i_clk 		=> clk,
		i_rst 		=> rst,
		i_speed		=> speed,
		o_current	=> c_base_pos,
		i_target	=> t_base_pos,
		o_pwm_out	=> b_pwm
	);


	movement 	: process(c_lower_pos, t_lower_pos, c_middle_pos, t_middle_pos, c_upper_pos, t_upper_pos)
	begin
		if((c_lower_pos = t_lower_pos) AND (c_middle_pos = t_middle_pos) AND (c_upper_pos = t_upper_pos)) then
			moving <= '0';
		else 
			moving <= '1';
		end if;

		l1 <= l_pwm;
		l2 <= l_pwm;
		m1 <= m_pwm;
		m2 <= m_pwm;
		u1 <= u_pwm;
		u2 <= u_pwm;
		g1 <= g_pwm;
		w1 <= w_pwm;
		b1 <= b_pwm;
		
	end process;
end v1;


